module rocketchip_wrapper (
    
)